module Sigmoid();
    
endmodule
