module sigmoid(x, z, clk);

	//Piecewise linear approximation

	input  signed [31:0] x;
	input  clk;
	output reg signed [31:0] y;
	
	wire signed [31:0] w1, w2;
	mult m1 (x, 0__0000_0100_0000_0000_0000_0000, w1);					//0.015625
	mult m2 (x, 0__0100_0000_0000_0000_0000_0000, w2);					//0.25

	
	always @(posedge clk)
	begin
		if (x + 1000__0000_0000_0000_0000_0000_0000 < 0)				//x + 8 < 0
			y <= 0;
			
		else if (x + 1__1001_1001_1001_1001_1001_1001 < 0)				//x + 1.6 < 0
			y <= 1000__0000_0000_0000_0000_0000_0000 + w1;				//z = 8 + x*0.015625
		
		else if (x - 1__1001_1001_1001_1001_1001_1001 < 0)				//x - 1.6 < 0
			y <= 0__1000_0000_0000_0000_0000_0000 + w2;					//z = 0.5 + x*0.25
		
		else if (x - 1000__0000_0000_0000_0000_0000_0000 < 0)			//x - 8 < 0
			y <= 0__1110_0000_0000_0000_0000_0000 - w1;					//z = 0.875 - x*0.015625
		
		else
			y <= 1__0000_0000_0000_0000_0000_0000;							//z = 1
	end

endmodule
